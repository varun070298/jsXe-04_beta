# JSXE Swedish properties file
# $Id: messages.sv,v 1.2 2006/02/16 21:29:20 ian_lewis Exp $
# Currently maintained by Patrik Johansson <patjoh@itstud.chalmers.se>
#:mode=properties:
#:tabSize=4:indentSize=4:noTabs=true:
#:folding=explicit:collapseFolds=1:

